/*
 * Avalon memory-mapped peripheral that generates VGA
 *
 * Stephen A. Edwards
 * Columbia University
 *
 * Register map:
 *
 * Byte Offset  7 ... 0   Meaning
 *        0    |  Red  |  Red component of background color (0-255)
 *        1    | Green |  Green component
 *        2    | Blue  |  Blue component
 *        3    | xlo   |  8 LSbs of the x-coordinate
 *        4    | xhi   |  3 MSbs of the x-coordinate (bits 7:3 are reserved)
 *        5    | ylo   |  8 LSbs of the y-coordinate
 *        6    | yhi   |  2 MSbs of the y-coordinate (bits 7:2 are reserved)
 */

`ifndef BALL_RADIUS_SQ
    `define BALL_RADIUS_SQ 21'h100 // 256
`endif
`ifndef BALL_INIT_X
    `define BALL_INIT_X 200
`endif
`ifndef BALL_INIT_Y
    `define BALL_INIT_Y 200
`endif

`define DRAW_BALL
`ifdef DRAW_BALL
module signed_mult_2_25(
    input  logic [26:0] a,
    input  logic [26:0] b,
    output logic [26:0] out);

    logic [53:0] mult_out;

    assign mult_out = a * b;
    assign out = mult_out[26:0];

endmodule
`endif

module vga_ball(input logic       clk,
                input logic       reset,
                input logic [7:0] writedata,
                input logic       write,
                input             chipselect,
                input logic [2:0] address,

                output logic [7:0] VGA_R, VGA_G, VGA_B,
                output logic       VGA_CLK, VGA_HS, VGA_VS,
                                   VGA_BLANK_n,
                output logic       VGA_SYNC_n);

    logic [10:0] hcount, next_hcount;
    logic [ 9:0] vcount;

    logic [ 7:0] background_r, background_g, background_b;
    logic [ 7:0] new_background_r, new_background_g, new_background_b;
    logic [10:0] ball_x;
    logic [10:0] new_ball_x;
    logic [ 9:0] ball_y;
    logic [ 9:0] new_ball_y;

`ifdef DRAW_BALL
    logic [10:0] dx, dx_q;
    logic [26:0] dx2;
    logic [ 9:0] dy, dy_q;
    logic [26:0] dy2;
    logic [21:0] dist2, dist2_q;
`endif

    vga_counters counters(.clk50(clk), .*);

`ifdef DRAW_BALL
    // calculate distance for the second future pixel
    // pipeline depth is 2 (1 pixel forward)
    assign next_hcount = hcount + 1;
    assign dx = (next_hcount >> 1) > ball_x ? (next_hcount >> 1) - ball_x : ball_x - (next_hcount >> 1);
    assign dy =      vcount > ball_y ?      vcount - ball_y : ball_y -      vcount;
    signed_mult_2_25 square_dx ( .a({16'b0, dx_q}), .b({16'b0, dx_q}), .out(dx2));
    signed_mult_2_25 square_dy ( .a({17'b0, dy_q}), .b({17'b0, dy_q}), .out(dy2));
    assign dist2 = dx2[21:0] + {2'b0, dy2[19:0]};

    always_ff @(posedge clk) begin
        if (reset) begin
            dx_q <= 11'b0;
            dy_q <= 10'b0;
            dist2_q <= 22'b0;
        end else begin
            dx_q <= dx;
            dy_q <= dy;
            dist2_q <= dist2;
        end
    end
`endif

    // take input from software
    always_ff @(posedge clk)
        if (reset) begin
            new_background_r <= 8'h0;
            new_background_g <= 8'h0;
            new_background_b <= 8'h80;
            new_ball_x       <= 11'd`BALL_INIT_X;
            new_ball_y       <= 10'd`BALL_INIT_Y;
        end else if (chipselect && write)
            case (address)
                3'h0 : new_background_r <= writedata;
                3'h1 : new_background_g <= writedata;
                3'h2 : new_background_b <= writedata;
                3'h3 : new_ball_x[ 7:0] <= writedata;
                3'h4 : new_ball_x[10:8] <= writedata[2:0];
                3'h5 : new_ball_y[ 7:0] <= writedata;
                3'h6 : new_ball_y[ 9:8] <= writedata[1:0];
            endcase

    // update control when starting a new frame (i.e., VGA_VS is high)
    always_ff @(posedge clk)
        if (reset) begin
            background_r <= 8'h0;
            background_g <= 8'h0;
            background_b <= 8'h80;
            ball_x       <= 11'd`BALL_INIT_X;
            ball_y       <= 10'd`BALL_INIT_Y;
        end else if (~VGA_VS) begin // new frame
        //end else begin
            background_r <= new_background_r;
            background_g <= new_background_g;
            background_b <= new_background_b;
            ball_x       <= new_ball_x;
            ball_y       <= new_ball_y;
        end

    // draw ball
    always_comb begin
        {VGA_R, VGA_G, VGA_B} = {8'h0, 8'h0, 8'h0};
        if (VGA_BLANK_n) begin
`ifdef DRAW_BALL
            // draw ball
            if (dist2_q < `BALL_RADIUS_SQ) begin
`else
            // draw rectangle in a box
            if (hcount[10:6] == ball_x[10:6] &&
                vcount[ 9:5] == ball_y[ 9:5]) begin
                {VGA_R, VGA_G, VGA_B} = {8'hff, 8'hff, 8'hff};
`endif
            end else begin
                {VGA_R, VGA_G, VGA_B} =
                    {background_r, background_g, background_b};
            end
        end
    end

endmodule

module vga_counters(
 input logic        clk50, reset,
 output logic [10:0] hcount,  // hcount[10:1] is pixel column
 output logic [9:0]  vcount,  // vcount[9:0] is pixel row
 output logic       VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n, VGA_SYNC_n);

/*
 * 640 X 480 VGA timing for a 50 MHz clock: one pixel every other cycle
 *
 * HCOUNT 1599 0             1279       1599 0
 *             _______________              ________
 * ___________|    Video      |____________|  Video
 *
 *
 * |SYNC| BP |<-- HACTIVE -->|FP|SYNC| BP |<-- HACTIVE
 *       _______________________      _____________
 * |____|       VGA_HS          |____|
 */
   // Parameters for hcount
   parameter HACTIVE      = 11'd 1280,
             HFRONT_PORCH = 11'd 32,
             HSYNC        = 11'd 192,
             HBACK_PORCH  = 11'd 96,
             HTOTAL       = HACTIVE + HFRONT_PORCH + HSYNC +
                            HBACK_PORCH; // 1600

   // Parameters for vcount
   parameter VACTIVE      = 10'd 480,
             VFRONT_PORCH = 10'd 10,
             VSYNC        = 10'd 2,
             VBACK_PORCH  = 10'd 33,
             VTOTAL       = VACTIVE + VFRONT_PORCH + VSYNC +
                            VBACK_PORCH; // 525

   logic endOfLine;

   always_ff @(posedge clk50 or posedge reset)
     if (reset)          hcount <= 0;
     else if (endOfLine) hcount <= 0;
     else            hcount <= hcount + 11'd 1;

   assign endOfLine = hcount == HTOTAL - 1;

   logic endOfField;

   always_ff @(posedge clk50 or posedge reset)
     if (reset)          vcount <= 0;
     else if (endOfLine)
       if (endOfField)   vcount <= 0;
       else              vcount <= vcount + 10'd 1;

   assign endOfField = vcount == VTOTAL - 1;

   // Horizontal sync: from 0x520 to 0x5DF (0x57F)
   // 101 0010 0000 to 101 1101 1111
   assign VGA_HS = !( (hcount[10:8] == 3'b101) &
            !(hcount[7:5] == 3'b111));
   assign VGA_VS = !( vcount[9:1] == (VACTIVE + VFRONT_PORCH) / 2);

   assign VGA_SYNC_n = 1'b0; // For putting sync on the green signal; unused

   // Horizontal active: 0 to 1279     Vertical active: 0 to 479
   // 101 0000 0000  1280         01 1110 0000  480
   // 110 0011 1111  1599         10 0000 1100  524
   assign VGA_BLANK_n = !( hcount[10] & (hcount[9] | hcount[8]) ) &
         !( vcount[9] | (vcount[8:5] == 4'b1111) );

   /* VGA_CLK is 25 MHz
    *             __    __    __
    * clk50    __|  |__|  |__|
    *
    *             _____       __
    * hcount[0]__|     |_____|
    */
   assign VGA_CLK = hcount[0]; // 25 MHz clock: rising edge sensitive

endmodule
