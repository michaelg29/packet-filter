
`include "packet_filter.svh"
`include "filter_defs.svh"

// Integrate input_fsm, type_field_checker, and dest_calculator
`timescale 1 ps / 1 ps
module preliminary_processor #(

) (
    input  logic clk,
    input  logic reset

);



endmodule
