
`include "packet_filter.svh"
`include "filter_defs.svh"

// Integrate sideband_buffer, frame_buffer, and switch_requester
`timescale 1 ps / 1 ps
module request_buffer #(

) (
    input  logic clk,
    input  logic reset

);



endmodule
