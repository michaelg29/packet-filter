
`ifndef _SYNTH_DEFS_SVH_
`define _SYNTH_DEFS_SVH_

`define TOP_TESTING
`define INTG_TESTING_1

`endif // _SYNTH_DEFS_SVH_
